`timescale 1ns / 1ps


module Mux_16x1_TB_v;

	// Inputs
	reg [15:0] I;
	reg [3:0] S;

	// Outputs
	wire O;

	// Instantiate the Unit Under Test (UUT)
	Mux_16x1 uut (
		.I(I), 
		.S(S), 
		.O(O)
	);

	initial begin
		// Initialize Inputs
		I = 0;
		S = 0;
		// Wait 100 ns for global reset to finish
		#5;
        
		I=16'b0000000000000001; S=4'b0000; #10;
		I=16'b0000000000000010; S=4'b0001; #10;
		I=16'b0000000000000100; S=4'b0010; #10;
		I=16'b0000000000001000; S=4'b0011; #10;
		I=16'b0000000000010000; S=4'b0100; #10;
		I=16'b0000000000100000; S=4'b0101; #10;
		I=16'b0000000001000000; S=4'b0110; #10;
		I=16'b0000000010000000; S=4'b0111; #10;
		I=16'b0000000100000000; S=4'b1000; #10;
		I=16'b0000001000000000; S=4'b1001; #10;
		I=16'b0000010000000000; S=4'b1010; #10;
		I=16'b0000100000000000; S=4'b1011; #10;
		I=16'b0001000000000000; S=4'b1100; #10;
		I=16'b0010000000000000; S=4'b1101; #10;
		I=16'b0100000000000000; S=4'b1110; #10;
		I=16'b1000000000000000; S=4'b1111; #10;
	end
endmodule

