`timescale 1ns / 1ps

module AND_GATE(A, B, F);
input A, B;
output F;

and(F, A, B);

endmodule
