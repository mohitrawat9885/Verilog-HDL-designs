`timescale 1ns / 1ps

module mohit_tb();
reg I0, I1, I2, I3, S0, S1;
wire Out;

mohit (I0, I1, I2, I3, S0, S1, Out);
initial
	begin
					 S1=0;S0=0;
					 I3=0;I2=0;I1=0;I0=0; #20;
					 I3=0;I2=0;I1=0;I0=1; #20;
					 I3=0;I2=0;I1=1;I0=0; #20;
					 I3=0;I2=0;I1=1;I0=1; #20;
				    I3=0;I2=1;I1=0;I0=0; #20;
					 I3=0;I2=1;I1=0;I0=1; #20;
					 I3=0;I2=1;I1=1;I0=0; #20;
					 I3=0;I2=1;I1=1;I0=1; #20;
					 
		          S1=0;S0=1;
					 I3=1;I2=0;I1=0;I0=0; #20;
					 I3=1;I2=0;I1=0;I0=1; #20;
					 I3=1;I2=0;I1=1;I0=0; #20;
					 I3=1;I2=0;I1=1;I0=1; #20;
				    I3=1;I2=1;I1=0;I0=0; #20;
					 I3=1;I2=1;I1=0;I0=1; #20;
					 I3=1;I2=1;I1=1;I0=0; #20;
					 I3=1;I2=1;I1=1;I0=1; #20;
		
				    S1=1;S0=0;
					 I3=0;I2=0;I1=0;I0=0; #20;
					 I3=0;I2=0;I1=0;I0=1; #20;
					 I3=0;I2=0;I1=1;I0=0; #20;
					 I3=0;I2=0;I1=1;I0=1; #20;
				    I3=0;I2=1;I1=0;I0=0; #20;
					 I3=0;I2=1;I1=0;I0=1; #20;
					 I3=0;I2=1;I1=1;I0=0; #20;
					 I3=0;I2=1;I1=1;I0=1; #20;
					 
					 S1=1;S0=1;
					 I3=1;I2=0;I1=0;I0=0; #20;
					 I3=1;I2=0;I1=0;I0=1; #20;
					 I3=1;I2=0;I1=1;I0=0; #20;
					 I3=1;I2=0;I1=1;I0=1; #20;
				    I3=1;I2=1;I1=0;I0=0; #20;
					 I3=1;I2=1;I1=0;I0=1; #20;
					 I3=1;I2=1;I1=1;I0=0; #20;
					 I3=1;I2=1;I1=1;I0=1; #20;
		
end
		
endmodule
