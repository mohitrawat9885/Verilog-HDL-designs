`timescale 1ns / 1ps

module NAND_GATE(A, F);
input A;
output F;

not(F, A);

endmodule
